** BJTOPT.SP BJT S-PARAMETER OPTIMIZATION
.OPTION ACCT NOMOD POST=2
* THE NET COMMAND IS AUTOMATICALLY REVERSING THE SIGN OF

* THE POWER SUPPLY CURRENT FOR THE NETWORK CALCULATIONS
.NET I(VCE) IBASE ROUT=50 RIN=50
VCE  VCE 0 10V
IBASE 0 IIN   AC=1 DC=.1MA
LBB  IIN BASE  #LBB#
LCC  VCE COLLECT #LCC#
LEE  EMIT 0 #LEE#

Q1 COLLECT BASE EMIT T2N6604
.MODEL T2N6604 NPN RB=#RB#  BF=100 TF=#TF# CJE=#CBE# CJC=#CBC#
+ RE=#RE# RC=#RC#  IS=#IS#

*.PARAM
*+ LBB= OPT1(100P, 1P, 10N)
*+ LCC= OPT1(100P, 1P, 10N)
*+ LEE= OPT1(100P, 1P, 10N)
*+ TF = OPT1(1N,  5P,  5N)
*+ CBE= OPT1(.5P, .1P, 5P)
*+ CBC= OPT1(.4P, .1P, 5P)
*+  RB= OPT1(10, 1, 300)
*+  RE= OPT1(.4, .01, 5)
*+  RC= OPT1(10, .1, 100)
*+  IS= OPT1(1E-15, 1E-16, 1E-10)
*.AC DATA=MEASURED  OPTIMIZE=OPT1
*+   RESULTS=COMP1,COMP3,COMP5,COMP6,COMP7
*+   MODEL=CONVERGE
.MODEL CONVERGE OPT RELIN=1E-4 RELOUT=1E-4 CLOSE=100 ITROPT=25
.MEASURE AC COMP1 ERR1 PAR(S11M) S11(M)
.MEASURE AC COMP2 ERR1 PAR(S11P) S11(P) MINVAL=10
.MEASURE AC COMP3 ERR1 PAR(S12M) S12(M)
.MEASURE AC COMP4 ERR1 PAR(S12P) S12(P) MINVAL=10
.MEASURE AC COMP5 ERR1 PAR(S21M) S21(M)
.MEASURE AC COMP6 ERR1 PAR(S21P) S21(P) MINVAL=10
.MEASURE AC COMP7 ERR1 PAR(S22M) S22(M)
.AC DATA=MEASURED
.PRINT PAR(S11M) S11(M) PAR(S11P) S11(P)
.PRINT PAR(S12M) S12(M) PAR(S12P) S12(P)
.PRINT PAR(S21M) S21(M) PAR(S21P) S21(P)
.PRINT PAR(S22M) S22(M) PAR(S22P) S22(P)
.DATA MEASURED
FREQ   S11M   S11P   S21M    S21P   S12M   S12P S22M   S22P
100ME  .6    -52     19.75   148    .02     65    .87   -21
200ME  .56   -95     15.30   127    .032    49    .69   -33
500ME  .56   -149     7.69    97    .044    41    .45   -41
1000ME .58   -174     4.07    77    .061    42    .39   -47
2000ME .61    159     2.03    50    .095    40    .39   -70
.ENDDATA
.PARAM FREQ=100ME S11M=0, S11P=0, S21M=0, S21P=0, S12M=0,
+  S12P=0, S22M=0, S22P=0
.END
.end





