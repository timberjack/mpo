*AMP.SP MOS OPERATIONAL AMPLIFIER OPTIMIZATION
.OPTION RELV=1E-3 RELVAR=.01 NOMOD ACCT POST
.PARAM VDD=5   VREF='VDD/2'
VDD VSUPPLY 0 VDD
VIN+    VIN+     0 PWL(0 ,'VREF-10M'   10NS 'VREF+10M' )
VINBAR+ VINBAR+  0 PWL(0 ,'VREF+10M'   10NS 'VREF-10M' )
VIN- VIN-  0  VREF
VBIAS VBIAS 0 #BIAS#
.GLOBAL VSUPPLY VBIAS

XRISE VIN+ VIN- VOUTR AMP
CLOADR VOUTR 0 .4P
XFALL VINBAR+ VIN- VOUTF AMP
CLOADF VOUTF 0 .4P

.MACRO AMP VIN+ VIN- VOUT
M1 2     VIN-   3       3       MOSN W=#WM1# L=#LM#
M2 4     VIN+   3       3       MOSN W=#WM1# L=#LM#
M3 2     2      VSUPPLY VSUPPLY MOSP W=#WM1# L=#LM#
M4 4     2      VSUPPLY VSUPPLY MOSP W=#WM1# L=#LM#
M5 VOUT  VBIAS  0       0       MOSN W=#WM5# L=#LM#
M6 VOUT  4      VSUPPLY VSUPPLY MOSP W=#WM6# L=#LM#
M7 3     VBIAS  0       0       MOSN W=#WM7# L=#LM#
.ENDS
.PARAM AREA='4*#WM1#*#LM# + #WM5#*#LM# + #WM6#*#LM# + #WM7#*#LM#'
VX 1000 0 AREA
RX 1000 0 1K
.MODEL MOSP PMOS (VTO=-1 KP=2.4E-5 LAMBDA=.004
+ GAMMA =.37 TOX=3E-8 LEVEL=3)
.MODEL MOSN NMOS (VTO=1.2 KP=6.0E-5 LAMBDA=.0004
+ GAMMA =.37 TOX=3E-8 LEVEL=3)

*.PARAM WM1=OPT1(60U,20U,100U)
*+      WM5=OPT1(40U,20U,100U)
*+      WM6=OPT1(300U,20U,500U)
*+      WM7=OPT1(70U,40U,200U)
*+       LM=OPT1(10U,2U,100U)
*+     BIAS=OPT1(2.2,1.2,3.0)

*.TRAN 2.5N 300N SWEEP OPTIMIZE=OPT1
*+     RESULTS=DELAYR,DELAYF,TOT_POWER,AREA_MIN  MODEL=OPT
*.MODEL OPT OPT CLOSE=100

.TRAN 2N 150N
.MEASURE DELAYR TRIG AT=0 TARG V(VOUTR) VAL=2.5 RISE=1
.MEASURE DELAYF TRIG AT=0 TARG V(VOUTF) VAL=2.5 FALL=1
.MEASURE TOT_POWER AVG POWER
.MEASURE AREA_MIN MIN PAR(AREA) MINVAL=100N
.PRINT V(VIN+) V(VOUTR) V(VOUTF)
.END
