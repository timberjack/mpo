*inverter based Oscillation Frequency
** HSPICE RF Simulation Options :
.option sim_accuracy=10		*simulation data accuracy
.option ingold=1			*science math. record (x.y*10ez)
.option POST=2				*control output ?
.option nomod				*not listing process file in data output file
.option filetype=ascii

.include "model013.lib_inc"
.include "/spice/vc_pwl.txt"

vdd vdd 0 1.2
vss vss 0 0
.load "/spice/vc_pwl.txt"
*vc vc 0 PWL ( 0.0u 0.05 0.1u 0.07 0.2u 0.12 0.3u 0.25 0.5u 0.36 0.6u 0.49 0.7u 0.61 0.8u 0.70 0.9u 0.73 1.1u 0.77 1.2u 0.88 1.6u 0.93 1.8u 1.1 )

.subckt vcdl_inv vdd vss out in v_c
mp out in vdd vdd pfet l=2u w=4u	$ name drain gate source bulk device length width
mn out in cn vss nfet l=1.6u w=1.6u
mc cn v_c vss vss nfet l=1.6u w=1.6u
.ends

*.subckt vcdl_inv vdd vss out in v_c
x1 vdd vss in1 in vc  vcdl_inv
x2 vdd vss in2 in1 vc  vcdl_inv
x3 vdd vss in3 in2 vc  vcdl_inv
x4 vdd vss in4 in3 vc  vcdl_inv
x5 vdd vss in5 in4 vc  vcdl_inv
x6 vdd vss in6 in5 vc  vcdl_inv
x7 vdd vss in7 in6 vc  vcdl_inv
x8 vdd vss in8 in7 vc  vcdl_inv
x9 vdd vss in9 in8 vc  vcdl_inv
x10 vdd vss in10 in9 vc  vcdl_inv
x11 vdd vss in11 in10 vc  vcdl_inv
x12 vdd vss in12 in11 vc  vcdl_inv
x13 vdd vss in13 in12 vc  vcdl_inv
x14 vdd vss in14 in13 vc  vcdl_inv
x15 vdd vss in15 in14 vc  vcdl_inv
x16 vdd vss in16 in15 vc  vcdl_inv
x17 vdd vss in17 in16 vc  vcdl_inv
x18 vdd vss in18 in17 vc  vcdl_inv
x19 vdd vss in in18 vc  vcdl_inv


*Transient Analysis Test Bench	$stimulate oscillation with 2mA pu
.ic v(in)=1.2 v(vc)=0.0
.tran 100p 10u

.save v(in) v(vc)
*.save @m.x3.mp[id]

*.control
*run
*set filetype=ascii
*write invo.txt v(in) v(vc)
*plot v(in) v(vc)
*plot (-1)*i(vdd)
*.endc

.END
