*Digital inverter

.PARAM V_SUPPLY = '3'
.PARAM INP_FREQ = '850000000'
.PARAM INP_PERIOD = '1/INP_FREQ'
.PARAM NO_PERIODS = '4'
.PARAM TMEAS_START = '(NO_PERIODS-1)*INP_PERIOD'
.PARAM TMEAS_STOP = '(NO_PERIODS)*INP_PERIOD'
.PARAM TMEAS_1 = 'TMEAS_STOP -3*INP_PERIOD/4'
.PARAM TMEAS_2 = 'TMEAS_STOP -1*INP_PERIOD/4'

*** *** SUPPLY VOLTAGES *** ***
VDD VDD 0 V_SUPPLY
VSS VSS 0 0

*** *** INPUT SIGNAL *** ***
VSIG IN VSS PULSE V_SUPPLY 0 'INP_PERIOD/2' 'INP_PERIOD/1000'
+               'INP_PERIOD/1000' 'INP_PERIOD/2' 'INP_PERIOD'

*** *** CIRCUIT *** ***
MP OUT IN VDD VDD PMOS W='0.005'   L=0.00001 pd='2*0.005+2*0.00000035' ps='2*0.005+2*0.00000035'
MN OUT IN VSS VSS NMOS W='0.005/3' L=0.00001 pd='2*0.005+2*0.00000035' ps='2*0.005+2*0.00000035'

CL OUT VSS 10p

*** *** ANALYSIS *** ***
.TRAN 'INP_PERIOD/1000' 'NO_PERIODS*INP_PERIOD'
*
*.PROBE TRAN V(IN)
.PROBE TRAN V(OUT)
.OPTION POST PROBE ACCURATE
.include p.typ
.include n.typ
.END

.measure tran P_SUPPLY rms par('i(vdd)*v_supply') from='tmeas_start' to='tmeas_stop'
.measure tran VHIGH find v(OUT) at='TMEAS_2'
.measure tran VLOW find v(OUT) at='TMEAS_1'

